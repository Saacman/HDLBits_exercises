module top_module (
    output out);
    assign out = 'b0;
endmodule